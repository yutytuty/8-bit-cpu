package types is
  type jmp_type_t is (T_JMP, T_JZ, T_JC, T_JS, T_JO, T_JA, T_JG, T_JGE);
end package;
